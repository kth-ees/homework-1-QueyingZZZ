`timescale 1ns/1ps

module arithmetic_right_shifter_tb;

  localparam N = 8;

  
  // complete
  // Inputs
endmodule
